library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 16;
          addrWidth: natural := 8
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  BEGIN
        -- Inicializa os endereços:
		  
tmp(0) := "0000101100000000";
tmp(1) := "0000110000001110";
tmp(2) := "0000100000000000";
tmp(3) := "0011011000001000";
tmp(4) := "0100001000000010";
tmp(5) := "0100001100000011";
tmp(6) := "0001010000000000";
tmp(7) := "0101000000001011";
tmp(8) := "0001010000000010";
tmp(9) := "0101000000001110";
tmp(10) := "0110000000010101";
tmp(11) := "0001010100000000";
tmp(12) := "0101000000010011";
tmp(13) := "0110000000010101";
tmp(14) := "0001010100000001";
tmp(15) := "0101000000010001";
tmp(16) := "0110000000010101";
tmp(17) := "0000101000001111";
tmp(18) := "0110000000010101";
tmp(19) := "0000101000001010";
tmp(20) := "0110000000010101";
tmp(21) := "0001011000000000";
tmp(22) := "0101000000011101";
tmp(23) := "0001011000000001";
tmp(24) := "0101000000011101";
tmp(25) := "0001011000000100";
tmp(26) := "0101000000100111";
tmp(27) := "0001011000000101";
tmp(28) := "0101000000100111";
tmp(29) := "0100010000000100";
tmp(30) := "0100010100000101";
tmp(31) := "0100000000000000";
tmp(32) := "0100000100000001";
tmp(33) := "0110000001000001";
tmp(34) := "0100010000000100";
tmp(35) := "0100010100000101";
tmp(36) := "0100110000000000";
tmp(37) := "0100101000000001";
tmp(38) := "0110000001000001";
tmp(39) := "0001101000001111";
tmp(40) := "0101000000101010";
tmp(41) := "0110000000100010";
tmp(42) := "0001010000000000";
tmp(43) := "0101000000101111";
tmp(44) := "0001010000000001";
tmp(45) := "0101000000101111";
tmp(46) := "0110000000111000";
tmp(47) := "1000010000001000";
tmp(48) := "0111010100000010";
tmp(49) := "0100010000000100";
tmp(50) := "0100010100000101";
tmp(51) := "0100110000000000";
tmp(52) := "0100101000000001";
tmp(53) := "0111010000001000";
tmp(54) := "1000010100000010";
tmp(55) := "0110000001000001";
tmp(56) := "0111010000000010";
tmp(57) := "0111010100000001";
tmp(58) := "0100010000000100";
tmp(59) := "0100010100000101";
tmp(60) := "0100110000000000";
tmp(61) := "0100101000000001";
tmp(62) := "1000010000000010";
tmp(63) := "1000010100000001";
tmp(64) := "0110000001000001";
tmp(65) := "0001011000000001";
tmp(66) := "0101000001110001";
tmp(67) := "0011100100000110";
tmp(68) := "0001100100000001";
tmp(69) := "0101000001000111";
tmp(70) := "0110000000000011";
tmp(71) := "0011100100000111";
tmp(72) := "0010000000000001";
tmp(73) := "0001000000001010";
tmp(74) := "0101000001001100";
tmp(75) := "0110000000000011";
tmp(76) := "0000000000000000";
tmp(77) := "0010000100000001";
tmp(78) := "0001000100000110";
tmp(79) := "0101000001010001";
tmp(80) := "0110000000000011";
tmp(81) := "0000000100000000";
tmp(82) := "0000100000000000";
tmp(83) := "0000100000000000";
tmp(84) := "0000100000000000";
tmp(85) := "0010001000000001";
tmp(86) := "0001001000001010";
tmp(87) := "0101000001011001";
tmp(88) := "0110000000000011";
tmp(89) := "0000001000000000";
tmp(90) := "0010001100000001";
tmp(91) := "0001001100000110";
tmp(92) := "0101000001011110";
tmp(93) := "0110000000000011";
tmp(94) := "0000001100000000";
tmp(95) := "0000100000000000";
tmp(96) := "0000100000000000";
tmp(97) := "0000100000000000";
tmp(98) := "0010010000000001";
tmp(99) := "0001010000001010";
tmp(100) := "0101000001101000";
tmp(101) := "0001010000000100";
tmp(102) := "0101000001101011";
tmp(103) := "0110000000000011";
tmp(104) := "0000010000000000";
tmp(105) := "0010010100000001";
tmp(106) := "0110000000000011";
tmp(107) := "0001010100000010";
tmp(108) := "0101000001101110";
tmp(109) := "0110000000000011";
tmp(110) := "0000010000000000";
tmp(111) := "0000010100000000";
tmp(112) := "0110000000000011";
tmp(113) := "0011011100001001";
tmp(114) := "0001011100000001";
tmp(115) := "0101000001110111";
tmp(116) := "0001011100000010";
tmp(117) := "0101000001111011";
tmp(118) := "0110000000000011";
tmp(119) := "0011011100001001";
tmp(120) := "0001011100000000";
tmp(121) := "0101000001010011";
tmp(122) := "0110000001110111";
tmp(123) := "0011011100001001";
tmp(124) := "0001011100000000";
tmp(125) := "0101000001100000";
tmp(126) := "0110000001111011";


--tmp(0) := "0011011000001000";
--tmp(1) := "0100000000000000";
--tmp(2) := "0100000100000001";
--tmp(3) := "0100001000000010";
--tmp(4) := "0100001100000011";
--tmp(5) := "0100010000000100";
--tmp(6) := "0100010100000101";
--tmp(7) := "0001011000000001";
--tmp(8) := "0101000000110111";
--tmp(9) := "0011100100000110";
--tmp(10) := "0001100100000001";
--tmp(11) := "0101000000001101";
--tmp(12) := "0110000000000000";
--tmp(13) := "0011100100000111";
--tmp(14) := "0010000000000001";
--tmp(15) := "0001000000001010";
--tmp(16) := "0101000000010010";
--tmp(17) := "0110000000000000";
--tmp(18) := "0000000000000000";
--tmp(19) := "0010000100000001";
--tmp(20) := "0001000100000110";
--tmp(21) := "0101000000010111";
--tmp(22) := "0110000000000000";
--tmp(23) := "0000000100000000";
--tmp(24) := "0000100000000000";
--tmp(25) := "0000100000000000";
--tmp(26) := "0000100000000000";
--tmp(27) := "0010001000000001";
--tmp(28) := "0001001000001010";
--tmp(29) := "0101000000011111";
--tmp(30) := "0110000000000000";
--tmp(31) := "0000001000000000";
--tmp(32) := "0010001100000001";
--tmp(33) := "0001001100000110";
--tmp(34) := "0101000000100100";
--tmp(35) := "0110000000000000";
--tmp(36) := "0000001100000000";
--tmp(37) := "0000100000000000";
--tmp(38) := "0000100000000000";
--tmp(39) := "0000100000000000";
--tmp(40) := "0010010000000001";
--tmp(41) := "0001010000001010";
--tmp(42) := "0101000000101110";
--tmp(43) := "0001010000000100";
--tmp(44) := "0101000000110001";
--tmp(45) := "0110000000000000";
--tmp(46) := "0000010000000000";
--tmp(47) := "0010010100000001";
--tmp(48) := "0110000000000000";
--tmp(49) := "0001010100000010";
--tmp(50) := "0101000000110100";
--tmp(51) := "0110000000000000";
--tmp(52) := "0000010000000000";
--tmp(53) := "0000010100000000";
--tmp(54) := "0110000000000000";
--tmp(55) := "0011011100001001";
--tmp(56) := "0001011100000001";
--tmp(57) := "0101000000111101";
--tmp(58) := "0001011100000010";
--tmp(59) := "0101000001000001";
--tmp(60) := "0110000000000000";
--tmp(61) := "0011011100001001";
--tmp(62) := "0001011100000000";
--tmp(63) := "0101000000011001";
--tmp(64) := "0110000000111101";
--tmp(65) := "0011011100001001";
--tmp(66) := "0001011100000000";
--tmp(67) := "0101000000100110";
--tmp(68) := "0110000001000001";




      return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 16;
          addrWidth: natural := 8
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  BEGIN
        -- Inicializa os endereços:
tmp(0) := "0011011000001000";
tmp(1) := "0100000000000000";
tmp(2) := "0100000100000001";
tmp(3) := "0100001000000010";
tmp(4) := "0100001100000011";
tmp(5) := "0100010000000100";
tmp(6) := "0100010100000101";
tmp(7) := "0001011000000001";
tmp(8) := "0101000000110111";
tmp(9) := "0011100100000110";
tmp(10) := "0001100100000001";
tmp(11) := "0101000000001101";
tmp(12) := "0110000000000000";
tmp(13) := "0011100100000111";
tmp(14) := "0010000000000001";
tmp(15) := "0001000000001010";
tmp(16) := "0101000000010010";
tmp(17) := "0110000000000000";
tmp(18) := "0000000000000000";
tmp(19) := "0010000100000001";
tmp(20) := "0001000100000110";
tmp(21) := "0101000000010111";
tmp(22) := "0110000000000000";
tmp(23) := "0000000100000000";
tmp(24) := "0000100000000000";
tmp(25) := "0000100000000000";
tmp(26) := "0000100000000000";
tmp(27) := "0010001000000001";
tmp(28) := "0001001000001010";
tmp(29) := "0101000000011111";
tmp(30) := "0110000000000000";
tmp(31) := "0000001000000000";
tmp(32) := "0010001100000001";
tmp(33) := "0001001100000110";
tmp(34) := "0101000000100100";
tmp(35) := "0110000000000000";
tmp(36) := "0000001100000000";
tmp(37) := "0000100000000000";
tmp(38) := "0000100000000000";
tmp(39) := "0000100000000000";
tmp(40) := "0010010000000001";
tmp(41) := "0001010000001010";
tmp(42) := "0101000000101110";
tmp(43) := "0001010000000100";
tmp(44) := "0101000000110001";
tmp(45) := "0110000000000000";
tmp(46) := "0000010000000000";
tmp(47) := "0010010100000001";
tmp(48) := "0110000000000000";
tmp(49) := "0001010100000010";
tmp(50) := "0101000000110100";
tmp(51) := "0110000000000000";
tmp(52) := "0000010000000000";
tmp(53) := "0000010100000000";
tmp(54) := "0110000000000000";
tmp(55) := "0011011100001001";
tmp(56) := "0001011100000001";
tmp(57) := "0101000000111101";
tmp(58) := "0001011100000010";
tmp(59) := "0101000001000001";
tmp(60) := "0110000000000000";
tmp(61) := "0011011100001001";
tmp(62) := "0001011100000000";
tmp(63) := "0101000000011001";
tmp(64) := "0110000000111101";
tmp(65) := "0011011100001001";
tmp(66) := "0001011100000000";
tmp(67) := "0101000000100110";
tmp(68) := "0110000001000001";




      return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;